
typedef enum bit {W, R} i2c_op_t;

